module camera_tb();

endmodule
