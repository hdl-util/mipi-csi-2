module camera_tb();
initial
begin
    $finish;
end
endmodule
